//Generating two 480 time-steps of 680 PRNG modules, storing them in an SRAM chip and displays them on a monitor via VGA protocol.
module High_arch_PRNG_VGA_SRAM(i_rst,SRAM_slot,i_clk,                                                //General declerations
i_CS_n,i_wr_trigger,i_rd_trigger,i_LB_n,i_UB_n,o_CS_n,o_OE_n,o_WE_n,o_LB_n,o_UB_n,o_A,I_O_bidir,     //SRAM declerations
o_red,o_green,o_blue,hsync,vsync,VGA_blank_N,VGA_sync_N,clk_25);                                     //VGA declerations
//Parameters
//PRNG parameters
parameter ARRAY_WIDTH=637;                             //Width of the one-dimensional CA grid
parameter i_arr_initial_value={318'd0,1'b1,318'd0};    //Initial value of the one-dimensional grid
parameter NEIGHBORHOOD=2;                              //Number of neuighboring cells
parameter N=10;                                        //Random number width. Not used in this TB.
parameter LOCATION=ARRAY_WIDTH/2;                      //Bit location for random number generation (input of the shift register). Not used in this TB.

//Input signals
input logic i_clk;                                     //50MHz clock
input logic i_rst;                                     //Active high logic. SW[0] in Altera DE2 board

input logic i_wr_trigger;                              //Trigerrs the write opration. Upon negative edge, 480 sequences of 640 bits are generated by the PRNG modules and stored in the SRAM memory. Key[0] in the DE-115 board.
input logic i_rd_trigger;                              //Trigerrs the read opration. Key[1] in the DE-115 board.
input logic SRAM_slot;                                 //When in Read mode, this switch chooses between upper- or lower-byte in the SRAM chip. SW[17] in Altera DE2 board.

input logic i_CS_n;                                    //SRAM chip select (active low). SW[1] in DE-115 board
input logic i_LB_n;                                    //SRAM lower-byte selection. SW[2] in DE-115 board.
input logic i_UB_n;                                    //SRAM upper-byte selection. SW[3] in DE-115 board.

//Output signals
//VGA output signals
output logic hsync;                                    //Horizontal sync signal
output logic vsync;                                    //Vertical sync signal
output logic [7:0]  o_red;                             //Input of the DAC in the VGA connector (converts into an analog signal between 0V-0.7V)
output logic [7:0]  o_green;                           //Input of the DAC in the VGA connector (converts into an analog signal between 0V-0.7V)
output logic [7:0]  o_blue;                            //Input of the DAC in the VGA connector (converts into an analog signal between 0V-0.7V)
output logic VGA_blank_N;                              //Tie to logic high (see ADV7123 video DAC datasheet)
output logic VGA_sync_N;                               //Tie to logic low (see ADV7123 video DAC datasheet)
output logic clk_25;                                   //25MHz clock


//SRAM output signals (SRAM cip IS61WV102416BLL)
output logic o_WE_n;                                   //SRAM write enable signal
output logic o_CS_n;                                   //SRAM chip-select signal
output logic o_LB_n;                                   //SRAM lower-byte enable signal
output logic o_UB_n;                                   //SRAM upper-byte enable signak
output logic o_OE_n;                                   //SRAM output enable (read) signal
output logic [19:0] o_A;                               //SRAM address bus

//SRAM data bus
inout logic [15:0] I_O_bidir;                          //SRAM data bus

//Internal signals
logic [ARRAY_WIDTH-1:0] o_sig_0;                       //Output word - m0 PRNG
logic [N-1:0] o_rn_0;                                  //N-bit random word
logic [ARRAY_WIDTH-1:0] o_sig_1;                       //Output word - m1 PRNG
logic [N-1:0] o_rn_1;                                  //N-bit random word

logic [9:0] count_n;                                   //SRAM controller internal counter, counts until ARRAY_WIDTH
logic [9:0] count_m;                                   //SRAM controller internal counter, count until 480
logic PRNG_en;                                         //Rises to logic high after the previous PRNG output has been written to the SRAM chip. Please see attached timing diagrams.
logic addr_inc;                                        //Rises to logic high when the VGA controller is at the 'active region'. It controls the address bus during read mode.

logic [15:0] I_O_tx;                                   //SRAM data bus - tx (bidir)
logic [15:0] I_O_rx;                                   //SRAM data bus - rx (bidir)

logic [9:0] next_x_cor;                                //X Coordinates of the next pixel
logic [9:0] next_y_cor;                                //y Coordinates of the next pixel

logic [7:0] i_color;                                   //VGA byte data
//HDL code

//25MHz clock generation
always @(posedge i_clk) 
  if (!i_rst)
    clk_25<=1'b0;
  else
    clk_25<=~clk_25;

//Instantiating CA_PRNG modules - Rule selection can be easialy modified via the 'RULE' parameter
CA_PRNG #(.ARRAY_WIDTH(ARRAY_WIDTH),.RULE(30),.NEIGHBORHOOD(NEIGHBORHOOD),.N(10),.LOCATION(LOCATION)) m0(.i_rst(i_rst),
                                                                                                         .i_clk(clk_25),
                                                                                                         .i_en(PRNG_en),
                                                                                                         .i_arr_initial_value(i_arr_initial_value),
                                                                                                         .o_sig(o_sig_0),
                                                                                                         .o_rn(o_rn_0)
);

CA_PRNG #(.ARRAY_WIDTH(ARRAY_WIDTH),.RULE(126),.NEIGHBORHOOD(NEIGHBORHOOD),.N(10),.LOCATION(LOCATION)) m1(.i_rst(i_rst),
                                                                                                         .i_clk(i_clk),
																																			.i_en(PRNG_en),
                                                                                                         .i_arr_initial_value(i_arr_initial_value),
                                                                                                         .o_sig(o_sig_1),
                                                                                                         .o_rn(o_rn_1)
);


//Instantiating N-bit to N-byte serial converters
//Upper byte
N_bit_to_N_Byte_converter #(.N(640), .COLOR_FORMAT(8'b11000100)) c1(.i_rst(i_rst&&~o_WE_n),
                                        .i_clk(clk_25),
                                        .i_data({{((640-ARRAY_WIDTH)/2){1'b0}},o_sig_0,{((640-ARRAY_WIDTH)/2+1){1'b0}}}), //Zero pedding the PRNG output sequence to 640
                                        .o_word(I_O_tx[15:8])
);
//Lower byte
N_bit_to_N_Byte_converter #(.N(640), .COLOR_FORMAT(8'b00101010)) c2(.i_rst(i_rst&&~o_WE_n),
                                        .i_clk(clk_25),
                                        .i_data({{((640-ARRAY_WIDTH)/2){1'b0}},o_sig_1,{((640-ARRAY_WIDTH)/2+1){1'b0}}}), //Zero pedding the PRNG output sequence to 640
                                        .o_word(I_O_tx[7:0])
);

//Instantiating SRAM controller (please see ocnceptual block and timing diagrams)
counter #(.N(640),.M(480)) c3(.i_rst(i_rst),
                              .i_clk(clk_25),
                              .i_en(o_WE_n),
                              .o_count_n(count_n),
                              .o_count_m(count_m)
);

control_signal_generator #(.N(640),.M(480)) c4(.i_rst(i_rst),
                                               .i_clk(clk_25),
                                               .i_count_n(count_n),
                                               .i_count_m(count_m),
                                               .i_wr_trigger(i_wr_trigger),
															  .i_rd_trigger(i_rd_trigger),
                                               .o_WE_n(o_WE_n),
															  .o_OE_n(o_OE_n),
                                               .o_PRNG_en(PRNG_en),
															  .i_next_x_cor(next_x_cor),
															  .i_next_y_cor(next_y_cor),
															  .o_addr_inc(addr_inc)
															  
);


address_counter #(.CNT_WIDTH(20)) c5 (.i_rst(i_rst),
                                      .i_wr_n(o_WE_n),
												  .i_rd_n(o_OE_n),
                                      .i_clk(clk_25),
												  .i_addr_inc(addr_inc),
                                      .A(o_A)
);

//SRAM data bus (bidir)
assign I_O_bidir = (o_WE_n==1'b1) ? 16'bzzzzzzzzzzzzzzzz : I_O_tx;
assign I_O_rx = I_O_bidir;

assign o_CS_n = i_CS_n;                                    //SRAM chip select signal
assign o_LB_n = i_LB_n;                                    //SRAM chip lower-byte enable signal
assign o_UB_n = i_UB_n;                                    //SRAM chip upper-byte enable signal

assign i_color = (SRAM_slot) ? (I_O_rx[7:0]) : (I_O_rx[15:8]);

//Instantiating the VGA driver
VGA_Driver v1(.i_rst(~o_OE_n),
              .i_clk(clk_25),
              .i_color(i_color),
              .hsync(hsync),
              .vsync(vsync),
              .o_red(o_red),
              .o_blue(o_blue),
              .o_green(o_green),
              .next_x_cor(next_x_cor),
              .next_y_cor(next_y_cor)
             );

assign VGA_blank_N=1'b1;                              //Tie to logic high (see ADV7123 video DAC datasheet)
assign VGA_sync_N=1'b0;                               //Tie to logic low (see ADV7123 video DAC datasheet)

endmodule
